module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
wire x,y,z,n;
    assign y= p2a&p2b;
    assign x= p2c&p2d;
    assign p2y= y|x;
    and(z,p1a,p1c,p1b);
    and(n,p1f,p1e,p1d);
    assign p1y= z|n;

endmodule
